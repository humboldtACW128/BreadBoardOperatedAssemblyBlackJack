PK   ���TւR`(  q�    cirkitFile.json��r$���_�A��H���\���9�X����{1Rt�
��0E��p,{z��2�6�=Ұ���E�Kτ}��L�~�����*$~��K+7����l�V��]��\�&y�]��?����//�^�l�o7�ޥ��]����]���mQ�]Iy��6����&�)���RNY�4�s	�{�6z�/^������ۂ�P7C��1����v3�Z����kAo|7C��	���f�f赠7c7C�����8G�'�nLH������e�	��O��&��?anMte}}�y���S���nLџu�M0��܇���:/"�^�齈>~�|�et�\�L�c��"B�E��zo������>�A���>��r�&�.��y���ﱻM0E��m�)���nL���v�`�~��m�)��N�	�F��S}�vX�y�b��S�g�?�;u����ߋ����twu�n�����i*�<U���i�ۄn��n
��������6�C��J�b�{�nL�ߣt���ߣt��MtS�*ӫD\�����WJ��N�ۄnb���w��Q�E��A�&����6��R��S�'�nLџ��Ml'"��M�w��������6���te�H�v�џ��MlgU�\iz��=�=9�Ey���ו}"�t^D��mb;E����&������N�	�	�z��S���&��_0,L<]�Lc�ݔo;����t�qc}GX�A�K�9�;�����tzc���X�A�K���;�����t<����c}�#,��X���t��ӛ��;(a��f��n��JGX:��X�E��t��k_f��`e��#0_���?��@��� �� ������}��Xe`���V ��VX>��`������|m��`Ł�#0_[p�Xu`������VX>��`������|�M0x��?�|�k����,���;_���o8Я8��À���,���z*�����G`���?�������a��?�|�k�����,��ںA�����G`����?�����o�>��B��a�#�|��U��od���G`�p`������|m5.�菴�_i����/X>��`������|�U˝����}�����p� ��V?X>�5�`������|mu>�`���#0_�+����,��ZE�����G`�V��?�|����Ձ �,_�|�k,��C�3A/4��/,_�|�ke?���,��Z������G`�Vj�?���������?�|�k�m���`���#0_���X`���j���X>�rD`������|���`���#0_���z�;z�;Xx���`���#0_+|�X`���Jv���X>�ja`������|����?�|�k����,��Zm9�����Gg������ޔ��M�a��*���MSR��b�\���|���+~l�ǚ��Y�T�rcqj�CR>TW�����W5�<�aA�'6?,��y(�����X�sn{�
��q�z�-���?~�!$3F\�j�'�ʺZ��^�O�}M�γ?��U���8�a�#�.�A��a
!+�C�S(�����k_���kg:Gn��1�s�<���A%��~暌	'ξ���g�>��2NvPN����*v6�C'U꾯j����i�<W�h�|������OA9�hO>﫚?~v[(U�-c���*�ɩ�svD5���8��揟�5NT�M�Ev]�CU��:̜ȋ=u����u�J5ƪ���[�L��ٍ��t*Ӯi��ٵO�4���Ю�H�(?�a�L�Z�:��揟�d����c�ǔ�K1���֖4�y>q�U�Oļ��f?�Z_�h����Tp%�1'�I�T̯i���S�6���r�G��8Uk�)��N�}U�γ?��W5<�s7�1�QFn�&�è�dl4��i8u��������vVs����R�Y�::�:&�ܔ���O�2F�ֆY��������9g�<�u��p*Ӯj�=�O������|{}{w��Ǐ���]0]�Vo�wq�|C�2��b�@�t{^0D C�=�"�!�q("�!��("�!��("�!�PD Cz3��@��&��@�Z!JX��em\چ�m�%n��V����K�?[k�;�`�e���1�28�R8��vc�f��C',��6�F�z�:���f3αv�+?d�!O�s`	��f�}Cb����K�.�N��7��t2m-��f���A�����M̝L�<����������Q�v[݃�`y���(Kz��=�	6����ϖ��O6GY��x��/�0�fRpS)���q���~� &�?YXGY�mV�qX��<����|�����Q�vӃ�`�q�Wq���q���&� &����Q�v;ă�`y����(K���AL�<�`yei��<f�����q��ݶ�91�{XGY��	���󸷛�כ�<�j�����q���n��L����Q�v[��^���x��q���6� �G,=�s���p��o�V�[�í�X��í�*������ p�@�J�.w��x�p�:�*Я����18\��
���rgy�W�í�*���u����p�@�J�.w��x�p<�*Я����18\�
���r'{�W�í�*����4��\�=�Acx�%B�����"}+$�dt�bz�Y�oe���^nP�7�����������f����`"�z��=�,ҷ22L�V/7�ǛE�VF����쑾�Qc"�$C��6�G�VF��В�����[U&BK2�m��̋]&BK2�m���oet�-�ж5W2�z#&�JLF�]fdt�-�ж5p2���e"�$C�����VF��Вm[�(�[]&BK2�mm��oet�-�ж5�2���e"�$C�ֺ��VF��Вm[���].��3��2IF��ж��2}��2Z��mk�e|+��DhI������׊B�+��2+�ˬ�.�%ڶ6_Ʒ2�L��dh[��q��.;B�6����.�2�L��dh[����2Z��m�+d|+��DhI������e"�$C�j���VF��Вm��"�[]&BK2�����oet�-�ж52�ZI&��LF�9]�dt�-�ж�A2���e"�$C�j��VF��Вm��$�[]&BK2����oet�-�ж�Z"��2�L��dh[m0���2Z��m5�d|+��DhI���j��.�%�VsNƷ2�L��dh[�<�
U�*�!�˼�.�2�L��dh[-C���2Z��m5e|+��DhI��Ֆ��.�%�V#SķAF��Вm��)�[]&BK2��f��oet�-��}�?6S��U�eVn����d�<����G7t~��Gj�>؟���L�UH5)7��9$��@uh{�Ws�e��#�m�h呚���b�N1���U9�7ݫ��笧��b�_BHf(|_�r�j5N��u�&�.9�`Yc�r���r��sF=�w�q�x~NC���P�J0,���e���~adGn��1�s�<���A%�8 rMƄ�,���e�>�l NvPN����*v6�#/U�"^VY9��"�jES�;m4[!��~
z�)F�&���r��FÆJU|�ٻ�LE79�}Ύ��0��,���eqC�ըFC�r���P�)�3�4Ů��UV���L�c�X?��*R��ϳ�/&�iE���Y�S M��-��2R)�y&��+XVY9�R��^������{5�b�s�-iN�|�e���ϑ��f?�Z_�h����Tp%�1'˽̊�h���,)g]��F�|Eq�j�S�Ƙ���<�*+����*+g�#�����#�u?1�Q��h
��"vWY9��d|����_gx(�j�*����7yZ���r�o4z�6�j��G�%E��ȩ*�/�m�}�*+Y~ښ���n�ݧ�r��Ǐf��9C�)�����C���� 2��C�@���9����3!��"��"b��"қE2�7#�dHo"�d�U=��H\�ƥmX�&X�FYj�iaL��M�䍲Ԫ�`��`	e�U߄1�r8��8�R��c��q��(K�� �	7���ay���8�R�c��q��(K���	��,��,�*W0&X7�<��Ԫ*��8,�[XGYjU|`L���T
,�[XGYj�V`L�<naye�U��1���q��VM�����Q�Z�,�;XGYj��aL�9qܤ8,�;XGYj��aL�<�`ye����1���q���j����=,��,�U�0&X��<���V���po7q�7ay���8�R[=c��q��(Km�
�	��,��,��0&X�<�����tX��A[�-H X%Va՛�*�U�_%XI�Uo+h�V�~�`%V�YT5@[�U��DXYw��uQ� �	Va�q��_� �`%V���uQ� �	Va՛E�U�_%XI�Uo�V�~�`%V�YT/@[�U��DX�7�2�@Fq�Вm��YƷB�KHv��.�^$��DhI��}k.�[�%BK2��y��(0Z��m����VF��Вm[� �[%&BK2�m-��oeԘ-�ж5%2��Qd"�$C�����VF��Вm[�#�bAF��Вm[�$�[]&BK2�m͕�o�ވ	���eFF�]&BK2�m��oet�-�ж�|2���e"�$C��$��VF��Вm[[)�[]&BK2�m���oet�-�ж��2���e"�$C����|�$��DhI���=��.�%ڶ�ZƷ2�L��dh�Zp�
}�(����.�2����2Z��mk�e|+��DhI�����.�%�V+AƷ2�L��dh[����2Z��m�+d|+��DhI������e"�$C�j���VF��Вm��"�[]&BK2�����oet�-�ж52�ZI&��LF�9]�dt�-�ж�A2���e"�$C�j��VF��Вm��$�[]&BK2����oet�-�ж�Z"��2�L��dh[m0���2Z��m5�d|+��DhI���j��.�%�VsNƷ2�L��dh[�<�
U�*�!�˼�.�2�L��dh[-C���2Z��m5e|+��DhI��Ֆ��.�%�V#SķAF��Вm��)�[]&BK2��f��oet�-��}��6S��U�eVn����d�<����G7t~��Gj�~��M�d�B�I��85�!)�C����,��`X�l�D+���h%Ku�AMu��9���^�\�8g=��+g�B2C���j��V�q"���5��u�q�+���h����h��0ꑽ��'��sBV.�:�P�aqt�/����#;rä�ɞ��AMF*��k2&�gYe�,K��Pfq��r:h��T���y�����Y~)�U+�*�i��
��S�CN1�5�e���,46T��{���f*�ɩ�svD5���gYe�,�j��F5����ݨ��L1u���)vE쮲r>�f*����	��U�ʤ|��X}1�N+��5Vβh�ij�m����JQ~��0��^����Y�������<f��s��ӞKomIs���,����|�4�AՒ��FT�+��9Y�eV<Gk��eI9��"�7��le�+��WC��5�Φ�YVY����VY9�q�� �|����Y�1�jH�FS8�������(%㣝���:�C�TkV���G���ӊ�h���}�ѣ�aV��<R-)��GNU)O|�l+��VYy���%����7������*���5��?\ݕw���i.ysu���������7G*�/\swc�6mpT�(��L��}�wi�-����I� Ci:���i*$J��,nгv���iOc7��K@�������S��t��t��tƁ�D��,���#�}r���B��#�;8���ƃ���eC=^����3��B��}jW$���ԙP�{��N��εU%�#p��+��3���w��u���]��g�vW���K�t����7�������˟/v���L��g� D��! x~hK���Ї����X?:����1t4}��F`���}�����$(�� �B! �)Q@��Fj��b��3xj�#�)�~�@���%����#�3��,���=5��d��%�T�x��a�����2_�+��$���]I��Nϊ*佅�g�P�_7}����~��d�˲O}'^�|���"���vN ���#����1 �7�Lr�m�_��n�ݧ�r�����ֺ;���v��*_�����m_9o���M�VvRt��ۯ�;)�M��W���&���St�`)�O�mBoB?E�	��)�M���O�mBob?E�	�Z���o�9��?	�@�m0 ����MH�s4z���sȪ�6��W�m0 ���ؾ�^��Yrڙ�ŊK��A�1�C��K���� R��%V�f:b�z_�%e�$������ ���������d�~m�c  �@Z��v�p Һ��ml��� ��-`�l�d��Q���ml��,.�wb!f%��1�d�~mC ���, ���ؾ�[\Z���b���6ڎl @.v�\�o�������`B������m��� G�7:����m�- �\� �~m+  �:@��]	����\�������W����= ����~ ����7v�Wv���|��r���~�o|�3~��= 5��hU��|�8 rq��V����ѽ�ioW&���b�$��Oo��q� ����Oo��q� ����Oo;e��A���#0K���`u^/���|<� �o��U��b���� ���Yu^/���|z�ع
g�?,���f�;��X>���b*�=���|�k_|��h&$4a�Z�C�
���!�!���}%��!Z��		MؾpF��H���&l�c�}�V%`BB�O��>D+0!�	�g�h��	��Є�~��
LHh¶� �C�J����@OT�u
��Єm�ڇh�&$4a[X��!��	��	Z��N1h�&$4a[���!Z��		M���}��)`BB��Qh�u
��Єm]ڇh�&$4a[���!Z��		M��ӡ}��)`BB.��^��_�����l�u��olвLHh¶�C�l��-E����k/�l�h�bѲLHh¶P�C�l�pY�����>���U��-�F�%Zŀ		M�Vs�}�V1`BB���h�U��Єm=؇-[���&l �>D�0!�	[��ѲLHh�V[�C�l��Յ@��N�P-[Z�8�l���@��S���&l�C�>D�0!�	[���:LHh�V��C�N����Уu
��Є�:ڇh�&$4a���!Z��		M���}��)`BB�Jh�u
��Є��ڇ�5��E�h���:ţu
��Є��ڇh�&$4a+
��!Z��		M�*��}��)`BB��k`�N��U�C��S���&lU��>D�0!�#�o�{{Sn�7��)S��2+7MIMd��u\py�Ñ�%��~Q��c{>�L&�*����S���q�:�bt5�ο�}����~Q&�c�P,�)5ձ*���Vzr���[�u�?q�!$3��]�j�'�ʺZ��^�O�M�������'�?�i�����q�z~�B���P�J0,N\���'���aR�dϭ�&����ۚk2&�:���'�}2��i�제Z%;U�l,�P����_�����ѡ<W�h�|����ķ�OA9�hO?��ڟ8?��M���α����nr*��QMa��ο����ƉjT��I����z��S���{�'�oU�S�/S��X5���;{�"�I�<���bb�N��5�O�_�HS��
�ڏT��C�Ʉ����j��%;�5�o3?����X�iO����9���j*�}�4�AՒ�"FT�+��9Y��'�M��O9��"���Gn?0��T�1�pn;u�U�{�"��j"�s���Fn�&��è�dl4��j8�ڟ�����vVs��"R�Y�::�R&dg�'�?��=Zf5��㷒�J~�$��ė�V��������?]^|lw�۾�l�]��|�(�������]|sy�f�����E��o[�5㥽3�`=Ӛ��ޙ�t�{���{�t�{��n{�tG�7rE���`M��k�&C�{iEJ�k�&�5�c��W<��1���|Ѐ���'�ܷs�?���n�M~I��1岧=�K(ꄢ�튼9e:�L���;e{�:�����덩�}#ͱ���������b�=Fz	�p8B8t�X�|.��3.��^��MV�>;�L��8�H���\��@��H�S_����ݣ�A_y_�~��NS�n]��Mmc�/��i�����-2~2˟쇟��'��'�����/
~
˟�?˟�?�˟⇟��'���t��jR!]_oܘ��z���zw�������l�|��pѯ�|�_u���y�y�v;���Q��_�}?n�髻۷����l��;&I7sika��ʷ���I߷�?8���o��=�#�9Po��*.���������|�����zyqW�������;���L7�r�7��G��h����Z�������0p����#�ǣ~������}{uۤ�<_��?�W��c��������i�z�^���;�����r��?��|�n�|��>�܃t��2�:?p/z�r;r~/
�x�~�l����-\f��,S�J�2(߄W![�8�|b0�ۛ�m�J:���]q�������|]>����+��+½Ü�� ���fk��W����n�R����K����X������zwwu���[�~�x{���9ڕ}�틣����r���wW�1y4d�O7�k���ߕ�S�����_����G���������*�Ʋ�������sI�����dMU4ǉ����k�?��U�(��sw��w�� ���ȸ|c�������φ�a���kѽ�fɺ���=+_� ���ƽز��v��3��Q�e�=r�K�ɶ�r�n/ۺ�l�j.���v�Hz���aG����D�#������������g�_�ݦ̗Fk�+
q�����I�ʒ��m���9�i�T��9���ڪ�15To�˚;��0W��X��,�G�gָdc����a��a/�#>�q_�h��ա7xV��zF�=a]�,{����^���7|V��|f��gq�K�HE��O>�7zV��~f�踐�Ǣgq�K�E��]ת��=qX<ˣ^&(�������E؏{�_���s�(V}��f�b9�{���Fhd�㿖��pP�㫾{n�/a��8F����%ƍ�N5����1��=���㿎�q�B�/�W}���?�z4�1J�%�%�|e�᫾&f�y���p��|�T�|�o���A��Vf��Ì���7_lߤ���'-H�W���8|�5�r��weG���4��1�\�
������|)��h���0�.�ț��@b�a98|?m�����f /�_�?3�zHڵ�0�Cw�]��fM�]~�t�u�n|�������5�8�<�X���d]����}��%��ؠ/�W�\|f|�I���΅w[>p���[s����E1�v4��Я�������*���d)��!���~W��{q�����o��=�|oX&W���]������/W��䛸����g������__�V�����_� :��uu���kY��`��s^o�ݥ�tQ�{?)�����_���3�O����oo�n�J��m-����__��$�_���.�ڿ�~�����ܸ��C���j֕G�p���3.��槯/~���HY�:x"6x�`�D��1����<z����^y��k�gq����.7O<Fc����т��0�Ckn8i�4�0��8a�x��$x���� O?��_>��K�>>�`���1���q;<�(ҏ�h�gq����������§�L�\,Y�1�c	��pڛn'>G�G�Q|�A+ǽ2�4`C)��Bi�#�}�4ǻ����ÿ>%�Z٩�f�c��a%T+�"=�\�<߶�l?1t�8��P���<jpG�:8���FDc��u�h��ɛ�*<<n��va���+�ZvOǂgm'V�61���Xh�81��P��9L�	�s
���;j���G��h����V���Q��sv��<<�U���3��9� xG=�y�,:x��@���`�`�&x���q?�:j|���Y���.��������]��)�ӻ�_����ߧ�������w_��.蛟.~�oPK
   ���TւR`(  q�                  cirkitFile.jsonPK      =   �(    